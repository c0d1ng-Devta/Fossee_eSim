* C:\eSim-Workspace\ALU\ALU.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/16/21 01:19:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ Net-_U4-Pad5_ Net-_U4-Pad6_ Net-_U4-Pad7_ Net-_U4-Pad8_ ALU		
v1  A1 Net-_R1-Pad2_ DC		
v2  A0 Net-_R2-Pad2_ DC		
v3  Net-_U2-Pad~_ Net-_R3-Pad2_ DC		
v4  Net-_U6-Pad~_ Net-_R4-Pad2_ DC		
v5  Net-_U3-Pad~_ Net-_R5-Pad2_ DC		
v6  Net-_U7-Pad~_ Net-_R6-Pad2_ DC		
U8  A1 A0 Net-_U2-Pad~_ Net-_U6-Pad~_ Net-_U3-Pad~_ Net-_U7-Pad~_ Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ Net-_U4-Pad5_ Net-_U4-Pad6_ adc_bridge_6		
U9  Net-_U4-Pad7_ Net-_U4-Pad8_ Net-_U11-Pad~_ Net-_U10-Pad~_ dac_bridge_2		
R1  GND Net-_R1-Pad2_ 1k		
R2  GND Net-_R2-Pad2_ 1k		
R3  GND Net-_R3-Pad2_ 1k		
R4  GND Net-_R4-Pad2_ 1k		
R5  GND Net-_R5-Pad2_ 1k		
R6  GND Net-_R6-Pad2_ 1k		
U11  Net-_U11-Pad~_ plot_v1		
U10  Net-_U10-Pad~_ plot_v1		
U5  A0 plot_v1		
U1  A1 plot_v1		
U2  Net-_U2-Pad~_ plot_v1		
U6  Net-_U6-Pad~_ plot_v1		
U3  Net-_U3-Pad~_ plot_v1		
U7  Net-_U7-Pad~_ plot_v1		

.end
